


// This module takes care of the control signal generation of the convolution operation
// based on the conv instruction

/*
module conv_ctr(
    input wire clk,
    input wire rst,
    input wire [3:0] current_kernel_size,
    input wire [8:0] current_feature_size

    output wire [3:0] kernel_size,
    output wire [8:0] feature_size
);*/